library verilog;
use verilog.vl_types.all;
entity system_memory_vlg_vec_tst is
end system_memory_vlg_vec_tst;
