LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY data_mem IS
	PORT(
		clk, wen, en	:	IN		STD_LOGIC;
		addr				:	IN		UNSIGNED(7 DOWNTO 0);
		data_in			:	IN 	STD_LOGIC_VECTOR(31 DOWNTO 0);
		data_out			:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
END data_mem;

ARCHITECTURE Behaviour OF data_mem IS

	TYPE RAM IS ARRAY (0 to 255) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL mem	:	RAM;
	
BEGIN

	PROCESS (wen, en, clk)
		BEGIN
			IF (clk' event AND clk = '0') THEN
				-- N/A
				IF	en = '0' THEN
					data_out <= (others => '0');
				-- read request
				ELSE
					IF wen = '0' THEN
						data_out <= mem(to_integer(addr));
					END IF;
				-- write request
					IF wen = '1' THEN
						mem(to_integer(addr)) <= data_in;
						data_out <= (others => '0');
					END IF;
				END IF;
			END IF;
	END PROCESS;
END Behaviour;